module memory(
    input clock, write_enable,
    input [31:0] address, data_in,
    output [31:0] data_out
);

endmodule